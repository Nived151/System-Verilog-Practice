//parameter